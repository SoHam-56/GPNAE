module PE5B (
    input wire [31:0] in,
    output reg [4:0] out
);
    always @(*) begin
        casez (in)
            32'b???????????????????????????????1: out = 5'd0;
            32'b??????????????????????????????10: out = 5'd1;
            32'b?????????????????????????????100: out = 5'd2;
            32'b????????????????????????????1000: out = 5'd3;
            32'b???????????????????????????10000: out = 5'd4;
            32'b??????????????????????????100000: out = 5'd5;
            32'b?????????????????????????1000000: out = 5'd6;
            32'b????????????????????????10000000: out = 5'd7;
            32'b???????????????????????100000000: out = 5'd8;
            32'b??????????????????????1000000000: out = 5'd9;
            32'b?????????????????????10000000000: out = 5'd10;
            32'b????????????????????100000000000: out = 5'd11;
            32'b???????????????????1000000000000: out = 5'd12;
            32'b??????????????????10000000000000: out = 5'd13;
            32'b?????????????????100000000000000: out = 5'd14;
            32'b????????????????1000000000000000: out = 5'd15;
            32'b???????????????10000000000000000: out = 5'd16;
            32'b??????????????100000000000000000: out = 5'd17;
            32'b?????????????1000000000000000000: out = 5'd18;
            32'b????????????10000000000000000000: out = 5'd19;
            32'b???????????100000000000000000000: out = 5'd20;
            32'b??????????1000000000000000000000: out = 5'd21;
            32'b?????????10000000000000000000000: out = 5'd22;
            32'b????????100000000000000000000000: out = 5'd23;
            32'b???????1000000000000000000000000: out = 5'd24;
            32'b??????10000000000000000000000000: out = 5'd25;
            32'b?????100000000000000000000000000: out = 5'd26;
            32'b????1000000000000000000000000000: out = 5'd27;
            32'b???10000000000000000000000000000: out = 5'd28;
            32'b??100000000000000000000000000000: out = 5'd29;
            32'b?1000000000000000000000000000000: out = 5'd30;
            32'b10000000000000000000000000000000: out = 5'd31;
            default: out = 5'b00000;
        endcase
    end
endmodule
